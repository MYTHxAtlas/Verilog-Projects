module inv_top_module(
	input in,
	output out);
	assign out = ~in;
endmodule
